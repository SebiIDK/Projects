** Profile: "SCHEMATIC1-R_cresc"  [ D:\Programe\Cadence\Laburi_Teme_Shit\Pop_Sebastian_Radu-PSpiceFiles\SCHEMATIC1\R_cresc.sim ] 

** Creating circuit file "R_cresc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../pop_sebastian_radu-pspicefiles/ledverde.lib" 
* From [PSPICE NETLIST] section of D:\Programe\Cadence\Working Shit\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM r 33k 66k 330 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
